module top_csi_fpga_wrapper_v #(
    localparam AXIM_ID_WIDTH     = 6,
    localparam AXIM_ADDR_WIDTH   = 48,
    localparam AXIM_DATA_WIDTH   = 32,
    localparam AXIM_USER_WIDTH   = 1,
    localparam AXIS_ID_WIDTH     = 1,
    localparam AXIS_ADDR_WIDTH   = 32,
    localparam AXIS_DATA_WIDTH   = 32,
    localparam AXIS_USER_WIDTH   = 1
)(
                    // clocks and reset interface
input wire                             reset_n_i,
input wire                             pixel_clk_i,
// AXI Slave Register Interface
input wire                              AXIS_ARESETN,
input wire                              AXIS_ACLK,
input           [AXIS_ADDR_WIDTH-1:0]   s_axi_awaddr,
input                                   s_axi_awvalid,
output wire                             s_axi_awready,

input           [AXIS_DATA_WIDTH-1:0]   s_axi_wdata,
input           [AXIS_DATA_WIDTH/8-1:0] s_axi_wstrb,
input                                   s_axi_wvalid,
output wire                             s_axi_wready,

output wire    [1:0]                    s_axi_bresp,
output wire                             s_axi_bvalid,
input                                   s_axi_bready,

input           [AXIS_ADDR_WIDTH-1:0]   s_axi_araddr,
input                                   s_axi_arvalid,
output  wire                            s_axi_arready,

output wire    [AXIS_DATA_WIDTH-1:0]    s_axi_rdata,
output wire    [1:0]                    s_axi_rresp,
output wire                             s_axi_rvalid,
input                                   s_axi_rready,

// AXI master interface
input wire                              AXIM_ACLK,
output wire    [AXIM_ID_WIDTH-1:0]      m_axi_awid,
output wire    [AXIM_ADDR_WIDTH-1:0]    m_axi_awaddr,
output wire    [7:0]                    m_axi_awlen,
output wire    [2:0]                    m_axi_awsize,
output wire    [1:0]                    m_axi_awburst,
output wire                             m_axi_awlock,
output wire    [3:0]                    m_axi_awcache,
output wire    [2:0]                    m_axi_awprot,
output wire    [3:0]                    m_axi_awqos,
output wire    [3:0]                    m_axi_awregion,
output wire    [5:0]                    m_axi_awatop,
//output wire    [AXIM_USER_WIDTH-1:0]    m_axi_awuser,
output wire                             m_axi_awvalid,
input                                   m_axi_awready,

output wire    [AXIM_DATA_WIDTH-1:0]    m_axi_wdata,
output wire    [AXIM_DATA_WIDTH/8-1:0]  m_axi_wstrb,
output wire                             m_axi_wlast,
//output wire    [AXIM_USER_WIDTH-1:0]    m_axi_wuser,
output wire                             m_axi_wvalid,
input                                   m_axi_wready,

input           [AXIM_ID_WIDTH-1:0]     m_axi_bid,
input           [1:0]                   m_axi_bresp,
//input           [AXIM_USER_WIDTH-1:0]   m_axi_buser,
input                                   m_axi_bvalid,
output wire                             m_axi_bready,

output wire    [AXIM_ID_WIDTH-1:0]      m_axi_arid,
output wire    [AXIM_ADDR_WIDTH-1:0]    m_axi_araddr,
output wire    [7:0]                    m_axi_arlen,
output wire    [2:0]                    m_axi_arsize,
output wire    [1:0]                    m_axi_arburst,
output wire                             m_axi_arlock,
output wire    [3:0]                    m_axi_arcache,
output wire    [2:0]                    m_axi_arprot,
output wire    [3:0]                    m_axi_arqos,
output wire    [3:0]                    m_axi_arregion,
//output wire    [AXIM_USER_WIDTH-1:0]    m_axi_aruser,
output wire                             m_axi_arvalid,
input  wire                             m_axi_arready,

input           [AXIM_ID_WIDTH-1:0]     m_axi_rid,
input           [AXIM_DATA_WIDTH-1:0]   m_axi_rdata,
input           [1:0]                   m_axi_rresp,
input                                   m_axi_rlast,
//input           [AXIM_USER_WIDTH-1:0]   m_axi_ruser,
input                                   m_axi_rvalid,
output wire                             m_axi_rready,
input wire                              rx_byte_clk_hs,
input wire                              rx_valid_hs0,
input wire                              rx_valid_hs1,
input wire                              rx_valid_hs2,
input wire                              rx_valid_hs3,
input wire      [7:0]                   rx_data_hs0,
input wire      [7:0]                   rx_data_hs1,
input wire      [7:0]                   rx_data_hs2,
input wire      [7:0]                   rx_data_hs3,
output wire                             frame_wr_done_intr
);
assign m_axi_awaddr[47:32] = 0;
assign m_axi_awid[5:1] = 0;
assign m_axi_arid[5:1] = 0;
top_csi_fpga_wrapper_sv top_csi_fpga_wrapper_sv_i(
    .reset_n_i              (   reset_n_i       ), 
    .pixel_clk_i            (   pixel_clk_i     ),

    // AXI Slave Interface
    .axi_clk_i              (   AXIS_ACLK       ),
    .axi_reset_n_i          (   AXIS_ARESETN    ),
    .s_axi_lite_awaddr_i    (   s_axi_awaddr    ),
    .s_axi_lite_awvalid_i   (   s_axi_awvalid   ),
    .s_axi_lite_awready_o   (   s_axi_awready   ),

    .s_axi_lite_wdata_i     (   s_axi_wdata     ),
    .s_axi_lite_wstrb_i     (   s_axi_wstrb     ),
    .s_axi_lite_wvalid_i    (   s_axi_wvalid    ),
    .s_axi_lite_wready_o    (   s_axi_wready    ),

    .s_axi_lite_bresp_o     (   s_axi_bresp     ),
    .s_axi_lite_bvalid_o    (   s_axi_bvalid    ),
    .s_axi_lite_bready_i    (   s_axi_bready    ),

    .s_axi_lite_araddr_i    (   s_axi_araddr    ),
    .s_axi_lite_arvalid_i   (   s_axi_arvalid   ),
    .s_axi_lite_arready_o   (   s_axi_arready   ),

    .s_axi_lite_rdata_o     (   s_axi_rdata     ),
    .s_axi_lite_rresp_o     (   s_axi_rresp     ),
    .s_axi_lite_rvalid_o    (   s_axi_rvalid    ),
    .s_axi_lite_rready_i    (   s_axi_rready    ),

    // AXI master interface
    .m_axi_csi_awid_o       (   m_axi_awid[0]      ),    
    .m_axi_csi_awaddr_o     (   m_axi_awaddr[31:0]    ),  
    .m_axi_csi_awlen_o      (   m_axi_awlen     ),   
    .m_axi_csi_awsize_o     (   m_axi_awsize    ),  
    .m_axi_csi_awburst_o    (   m_axi_awburst   ), 
    .m_axi_csi_awlock_o     (   m_axi_awlock    ),  
    .m_axi_csi_awcache_o    (   m_axi_awcache   ), 
    .m_axi_csi_awprot_o     (   m_axi_awprot    ),  
    .m_axi_csi_awqos_o      (   m_axi_awqos     ),   
    .m_axi_csi_awregion_o   (   m_axi_awregion  ),
    .m_axi_csi_awatop_o     (   m_axi_awatop    ),  
    .m_axi_csi_awuser_o     (   m_axi_awuser    ),  
    .m_axi_csi_awvalid_o    (   m_axi_awvalid   ), 
    .m_axi_csi_awready_i    (   m_axi_awready   ), 

    .m_axi_csi_wdata_o      (   m_axi_wdata     ),   
    .m_axi_csi_wstrb_o      (   m_axi_wstrb     ),   
    .m_axi_csi_wlast_o      (   m_axi_wlast     ),   
    .m_axi_csi_wuser_o      (   m_axi_wuser     ),   
    .m_axi_csi_wvalid_o     (   m_axi_wvalid    ),  
    .m_axi_csi_wready_i     (   m_axi_wready    ),  

    .m_axi_csi_bid_i        (   m_axi_bid[0]       ),     
    .m_axi_csi_bresp_i      (   m_axi_bresp     ),   
    .m_axi_csi_buser_i      (   m_axi_buser     ),   
    .m_axi_csi_bvalid_i     (   m_axi_bvalid    ),  
    .m_axi_csi_bready_o     (   m_axi_bready    ),  

    .m_axi_csi_arid_o       (   m_axi_arid[0]      ),    
    .m_axi_csi_araddr_o     (   m_axi_araddr[31:0]    ),  
    .m_axi_csi_arlen_o      (   m_axi_arlen     ),   
    .m_axi_csi_arsize_o     (   m_axi_arsize    ),  
    .m_axi_csi_arburst_o    (   m_axi_arburst   ), 
    .m_axi_csi_arlock_o     (   m_axi_arlock    ),  
    .m_axi_csi_arcache_o    (   m_axi_arcache   ), 
    .m_axi_csi_arprot_o     (   m_axi_arprot    ),  
    .m_axi_csi_arqos_o      (   m_axi_arqos     ),   
    .m_axi_csi_arregion_o   (   m_axi_arregion  ),
    .m_axi_csi_aruser_o     (   m_axi_aruser    ),
    .m_axi_csi_arvalid_o    (   m_axi_arvalid   ),
    .m_axi_csi_arready_i    (   m_axi_arready   ),

    .m_axi_csi_rid_i        (   m_axi_rid       ),
    .m_axi_csi_rdata_i      (   m_axi_rdata     ),
    .m_axi_csi_rresp_i      (   m_axi_rresp     ),
    .m_axi_csi_rlast_i      (   m_axi_rlast     ),
    .m_axi_csi_ruser_i      (   m_axi_ruser     ),
    .m_axi_csi_rvalid_i     (   m_axi_rvalid    ),
    .m_axi_csi_rready_o     (   m_axi_rready    ),
    .rx_byte_clk_hs_i       (   rx_byte_clk_hs  ),
    .rx_valid_hs0_i         (   rx_valid_hs0    ),
    .rx_valid_hs1_i         (   rx_valid_hs1    ),
    .rx_valid_hs2_i         (   rx_valid_hs2    ),
    .rx_valid_hs3_i         (   rx_valid_hs3    ),
    .rx_data_hs0_i          (   rx_data_hs0     ),
    .rx_data_hs1_i          (   rx_data_hs1     ),
    .rx_data_hs2_i          (   rx_data_hs2     ),
    .rx_data_hs3_i          (   rx_data_hs3     ),
    .frame_wr_done_intr_o   (frame_wr_done_intr )
);

endmodule
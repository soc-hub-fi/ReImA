module mem_write_axi(
                // input pixel interface
                input reset_n_i,
                input clk_i,
                input pixel_data_valid_i,
                input [63:0] pixel_data_i,
                // axi4 output interface
                output 
);

endmodule